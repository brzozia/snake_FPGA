library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity snake_vhdl is
port(
	reset, clk: in std_logic;
	a1,a2,b1,b2,c1,c2,d1,d2,e1,e2,f1,f2,g1,g2: out std_logic
	);
end snake_vhdl;



architecture arch1 of snake_vhdl is

--signal num: std_logic_vector(3 downto 0);	

variable num : integer;
begin

	process(num)

	begin
	
	
	case num is
		when 0 => 
			a1<='1';
			a2<='1';
			b2<='1';
			g2<='0';
			g1<='0';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';

			--(a1,a2,b2) <= ("1", "1","1");
			--(b1,c1,c2,d1,d2,e1,e2,f1,f2,g1,g2)<="00000000000";
			
		when 1 => 
			a1<='0';
			a2<='1';
			b2<='1';
			g2<='1';
			g1<='0';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
		
			--(a2, b2, g2}<=3'b111;
			--(b1,c1,c2,d1,d2,e1,e2,f1,f2,g1,a1)<=11'b00000000000;
			
		when 2 => 
			a1<='0';
			a2<='0';
			b2<='1';
			g2<='1';
			g1<='1';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(b2, g2, g1)<=3'b111;
			--(b1,c1,c2,d1,d2,e1,e2,f1,f2,a1,a2)<=11'b00000000000;
			
		when 3 => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='1';
			g1<='1';
			e1<='1';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(g2, g1, e1)<=3'b111;
			--(b1,c1,c2,d1,d2,e2,f1,f2,a1,a2,b2)<=11'b00000000000;
			
		when 4 => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='0';
			g1<='1';
			e1<='1';
			d1<='1';
			d2<='0';
			c2<='0';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(g1, e1,d1)<=3'b111;
			--(b1,c1,c2,d2,e2,f1,f2,a1,a2,b2,g2)<=11'b00000000000;
			
		when 5 => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='0';
			g1<='0';
			e1<='1';
			d1<='1';
			d2<='1';
			c2<='0';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(e1,d1,d2)<=3'b111;
			--(b1,c1,c2,e2,f1,f2,a1,a2,b2,g2,g1)<=11'b00000000000;
			
		when 6 => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='0';
			g1<='0';
			e1<='0';
			d1<='1';
			d2<='1';
			c2<='1';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
		--	(d1,d2,c2)<=3'b111;
--(b1,c1,e2,f1,f2,a1,a2,b2,g2,g1,e1)<=11'b00000000000;
			
		when 7 => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='1';
			g1<='0';
			e1<='0';
			d1<='0';
			d2<='1';
			c2<='1';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(d2,c2,g2)<=3'b111;
			--(b1,c1,e2,f1,f2,a1,a2,b2,g1,e1,d1)<=11'b00000000000;
			
		when 8 => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='1';
			g1<='1';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='1';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(c2,g2,g1)<=3'b111;
			--(b1,c1,e2,f1,f2,a1,a2,b2,e1,d1,d2)<=11'b00000000000;
			
		when 9 => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='1';
			g1<='1';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='1';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(g2,g1,f1)<=3'b111;
			--(b1,c1,e2,f2,a1,a2,b2,e1,d1,d2,c2)<=11'b00000000000;
			
		when 10 => 
			a1<='1';
			a2<='0';
			b2<='0';
			g2<='0';
			g1<='1';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='1';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(g1,f1,a1)<=3'b111;
			--(b1,c1,e2,f2,a2,b2,e1,d1,d2,c2,g2)<=11'b00000000000;
			
		when 11 => 
			a1<='1';
			a2<='1';
			b2<='0';
			g2<='0';
			g1<='0';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='1';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(f1,a1,a2)<=3'b111;
			--(b1,c1,e2,f2,b2,e1,d1,d2,c2,g2,g1)<=11'b00000000000;
			
		when others => 
			a1<='0';
			a2<='0';
			b2<='0';
			g2<='0';
			g1<='0';
			e1<='0';
			d1<='0';
			d2<='0';
			c2<='0';
			f1<='0';
			b1<='0';
			c1<='0';
			f2<='0';
			e2<='0';
			--(a1,a2,b1,b2,c1,c2,d1,d2,e1,e2,f1,f2,g1,g2)<=14'b00000000000000;
	
	end case;
end process;

	P2: process (clk)
	begin
		if rising_edge(clk) then
			if(reset='1')then num:=0;
			else
				if(num=11) then num:=0;
				else num:=num+1;
				end if;
			end if;
		end if;
	end process P2;
	
end arch1;




--case num is
--		when 0 => 
--			a1<='1';
--			a2<="1";
--			b2<="1";
--			g2<="0";
--			g1<="0";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			e2<="0";
--
--			--(a1,a2,b2) <= ("1", "1","1");
--			--(b1,c1,c2,d1,d2,e1,e2,f1,f2,g1,g2)<="00000000000";
--			
--		when 1 => 
--			a1<="0";
--			a2<="1";
--			b2<="1";
--			g2<="1";
--			g1<="0";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			e2<="0";
--		
--			--(a2, b2, g2}<=3'b111;
--			--(b1,c1,c2,d1,d2,e1,e2,f1,f2,g1,a1)<=11'b00000000000;
--			
--		when 2 => 
--			a1<="0";
--			a2<="0";
--			b2<="1";
--			g2<="1";
--			g1<="1";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			e2<="0";
--			--(b2, g2, g1)<=3'b111;
--			--(b1,c1,c2,d1,d2,e1,e2,f1,f2,a1,a2)<=11'b00000000000;
--			
--		when 3 => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="1";
--			g1<="1";
--			e1<="1";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(g2, g1, e1)<=3'b111;
--			--(b1,c1,c2,d1,d2,e2,f1,f2,a1,a2,b2)<=11'b00000000000;
--			
--		when 4 => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="0";
--			g1<="1";
--			e1<="1";
--			d1<="1";
--			d2<="0";
--			c2<="0";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(g1, e1,d1)<=3'b111;
--			--(b1,c1,c2,d2,e2,f1,f2,a1,a2,b2,g2)<=11'b00000000000;
--			
--		when 5 => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="0";
--			g1<="0";
--			e1<="1";
--			d1<="1";
--			d2<="1";
--			c2<="0";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(e1,d1,d2)<=3'b111;
--			--(b1,c1,c2,e2,f1,f2,a1,a2,b2,g2,g1)<=11'b00000000000;
--			
--		when 6 => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="0";
--			g1<="0";
--			e1<="0";
--			d1<="1";
--			d2<="1";
--			c2<="1";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--		--	(d1,d2,c2)<=3'b111;
----(b1,c1,e2,f1,f2,a1,a2,b2,g2,g1,e1)<=11'b00000000000;
--			
--		when 7 => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="1";
--			g1<="0";
--			e1<="0";
--			d1<="0";
--			d2<="1";
--			c2<="1";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(d2,c2,g2)<=3'b111;
--			--(b1,c1,e2,f1,f2,a1,a2,b2,g1,e1,d1)<=11'b00000000000;
--			
--		when 8 => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="1";
--			g1<="1";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="1";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(c2,g2,g1)<=3'b111;
--			--(b1,c1,e2,f1,f2,a1,a2,b2,e1,d1,d2)<=11'b00000000000;
--			
--		when 9 => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="1";
--			g1<="1";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="1";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(g2,g1,f1)<=3'b111;
--			--(b1,c1,e2,f2,a1,a2,b2,e1,d1,d2,c2)<=11'b00000000000;
--			
--		when 10 => 
--			a1<="1";
--			a2<="0";
--			b2<="0";
--			g2<="0";
--			g1<="1";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="1";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(g1,f1,a1)<=3'b111;
--			--(b1,c1,e2,f2,a2,b2,e1,d1,d2,c2,g2)<=11'b00000000000;
--			
--		when 11 => 
--			a1<="1";
--			a2<="1";
--			b2<="0";
--			g2<="0";
--			g1<="0";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="1";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(f1,a1,a2)<=3'b111;
--			--(b1,c1,e2,f2,b2,e1,d1,d2,c2,g2,g1)<=11'b00000000000;
--			
--		when others => 
--			a1<="0";
--			a2<="0";
--			b2<="0";
--			g2<="0";
--			g1<="0";
--			e1<="0";
--			d1<="0";
--			d2<="0";
--			c2<="0";
--			f1<="0";
--			b1<="0";
--			c1<="0";
--			f2<="0";
--			--(a1,a2,b1,b2,c1,c2,d1,d2,e1,e2,f1,f2,g1,g2)<=14'b00000000000000;
--	
--	end case;